module mux2(d0,d1,s,y);
input[31:0] d0, d1;	
input s;		
output [31:0] y;	
assign y = s ? d1 : d0 ;

endmodule

module mux3(d0,d1,d2,s,y);
input[31:0] d0, d1,d2;	
input[1:0] s;		
output reg [31:0] y;	
always @ (*)
begin
	case(s)
		2'b00:y = d0;
		2'b01:y = d1;
		2'b10:y = d2;
	endcase
end
endmodule

module mux4(d0,d1,d2,d3,s,y);
input[31:0] d0, d1,d2,d3;	
input[1:0] s;		
output reg [31:0] y;	
always @ (*)
begin
	case(s)
		2'b00:y = d0;
		2'b01:y = d1;
		2'b10:y = d2;
		2'b11:y = d3;
	endcase
end
endmodule
